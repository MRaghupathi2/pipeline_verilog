module pcadder(in,out);

input [15:0] in;
output [15:0] out;

assign out = in + 16'd1;

endmodule